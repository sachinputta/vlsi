module pri256_tb();
reg [255:0]d_in;
wire [255:0]d_out;
wire v;

pri256 pwe(d_out,d_in);

initial
begin
d_in=256'd01010101111100000000000000011101010101010000000000000;
#10
d_in=256'b000000000000000001111111111111110000000000001111111111110000;
#10
d_in=256'b01010101010101010101010100_0000_0000_0000_0000_0000_0000_0000_0000_0000;
end

initial
begin
$monitor($time," input=%b  pri_output=%b",d_in,d_out);
end
endmodule


module program(add,out);

input [4:0] add ;
output [31:0] out ;
reg [31:0] out ;


reg  [31:0]  PMEMORY [31:0];


always @(*) begin

        out = PMEMORY[add];
        
end

initial begin

PMEMORY[0]  = 32'b10000000010000000000000000000001;
PMEMORY[1]  = 32'b10000000100000000000000000000010;
PMEMORY[2]  = 32'b10000000110000000000000000000011;
PMEMORY[3]  = 32'b10000001000000000000000000000100;
PMEMORY[4]  = 32'b10000001010000000000000000000101;
PMEMORY[5]  = 32'b10000001100000000000000000000110;
PMEMORY[6]  = 32'b10000001110000000000000000000111;
PMEMORY[7]  = 32'b10000010000000000000000000001000;
PMEMORY[8]  = 32'b10000010010000000000000000001001;
PMEMORY[9]  = 32'b10000010100000000000000000001010;
PMEMORY[10] = 32'b10000010110000000000000000001011;
PMEMORY[11] = 32'b10000011000000000000000000001100;
PMEMORY[12] = 32'b10000011010000000000000000001101;
PMEMORY[13] = 32'b10000011100000000000000000001110;
PMEMORY[14] = 32'b10000011110000000000000000001111;
PMEMORY[15] = 32'b10000100000000000000000000010000;
PMEMORY[16] = 32'b10000100010000000000000000010001;
PMEMORY[17] = 32'b10000100100000000000000000010010;
PMEMORY[18] = 32'b
PMEMORY[19] = 32'b
PMEMORY[20] = 32'b
PMEMORY[21] = 32'b
PMEMORY[22] = 32'b
PMEMORY[23] = 32'b
PMEMORY[24] = 32'b
PMEMORY[25] = 32'b
PMEMORY[26] = 32'b





end

endmodule



module faddsub_tb();

reg [31:0]a,b;
reg clk;
wire [31:0]c;

fpa f1(a,b,c,clk);

initial 
begin

clk=1'b1;


a=32'b01101011111100111010000011000011;
b=32'b01101011100011100101111100011100;

#4
a=32'b00111111100110000000000000000000;
b=32'b00111111000100000000000000000000;
/*
#4

a=32'b00000000110100011110110000100000;
b=32'b00000000011001010001111011000010;
#4

a=32'b00000000110100011110110000100000;
b=32'b00000000011001010001111011000010;

#4

a=32'b00000000110100011110110000100000;
b=32'b00000000011001010001111011000010;


#4
a=32'b00000000110100011110110000100000;
b=32'b00000000011001010001111011000010;

#4
a=32'b00000000110100011110110000100000;
b=32'b00000000011001010001111011000010;*/

#32 $finish;
end

always
#2 clk=~clk;
initial
begin
$monitor("a=%b,b=%b,c=%b\n",a,b,c);
end
endmodule









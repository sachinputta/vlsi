      	 module ALU_tb();

reg [31:0]a2,a3,a4,a5,a6;
reg [31:0]b2,b3,b4,b5,b6,term1,term2;
reg [63:0]term3,term4,term5,term6,term7;
//reg [4:0]opcode;
wire [63:0]OUT,L11,L12,L13,L21,L22;


//tan18
//taylor series till first 7 terms\


//level 1
ALU l11(term1,term2,0101,L11);
ALU l12(term3[31:0],term4[31:0],0101,L12);
ALU l13(term5[31:0],term6[31:0],0101,L13);

//level 2
ALU l21(L11[31:0],L12[31:0],0101,L21);
ALU l22(term7[31:0],L13[31:0],0101,L22);	

//level 3
ALU l31(L21[31:0],L22[31:0],0101,OUT);

initial
begin
	term1=32'b01000001100010010000000000000000; 	        //18
	term2=32'b01000100100000111100110000000000;		//1944.00
	term3=32'b01001000011110110000010011001100;		//251942.4
	term4=32'b010010111111111000001010000011111;		//33040446.171428571
	term5=32'b010011111101000111111110101100011;		//5502584341.3046
	term6=32'b010100101111111011011110010011100;		//544895546735.57610
	term7=32'b010101101100010000001000110010010;		//74804530933100.67
end	

initial	
begin
$monitor(“tan(18)=%b\n”,OUT[31:0]);
end 	

endmodule // ALU_tb


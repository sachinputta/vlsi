module mresult_normalize(Mc,Sc,Ec,ScOut,EcOut,Mc1);
input [48:0]Mc;
input [7:0]Ec;
input Sc;
reg [48:0]McOut;
output reg [24:0]Mc1;
output reg [7:0]EcOut;
output reg ScOut;
always@ (*)
begin
     
     McOut= Mc;
     ScOut=Sc;
     EcOut=Ec; 
     Mc1[24:0]=McOut[48:24];
     $display("\nMc1[24]=%b\n",Mc1[24]);
	if(Mc1[24]==1'b1)
	begin
		Mc1=Mc1>>1'b1;
		EcOut=EcOut+8'b00000001;
		//$display("\nEntered if condition in result result_normalize now the McOut is %b\n",Mc1);
	end
	else
	begin
		
		repeat(24)
		begin
			if(Mc1[23]==1'b0)
			begin
				Mc1= Mc1<<1'b1;
				EcOut=EcOut-8'b00000001;
				//$display("\nEntered else condition in result result_normalize now the McOut is %b and EcOut is %b\n",Mc1,EcOut);
			end
		end	
	end
	
end

	
	

endmodule

module mcarry_calculation(a,b,p,cin,c);
  input [47:0]a,b;
  input cin;
  output [47:0]p;
  wire [47:0]g;
  output [48:0]c;  
  
assign g=a&b;

assign p=a^b;
  
assign c[0]=g[0]|(p[0]&cin);

assign c[1]=g[1]|(p[1]&(g[0]|(p[0]&cin)));

assign c[2]=g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))));

assign c[3]=g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))));

assign c[4]=g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))));

assign c[5]=g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))));

assign c[6]=g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))));

assign c[7]=g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))));

assign c[8]=g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))));

assign c[9]=g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))));

assign c[10]=g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))));

assign c[11]=g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))));

assign c[12]=g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))));

assign c[13]=g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))));

assign c[14]=g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))));

assign c[15]=g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))));

assign c[16]=g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))));

assign c[17]=g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))));

assign c[18]=g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))));

assign c[19]=g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))));

assign c[20]=g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))));

assign c[21]=g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))));

assign c[22]=g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))));

assign c[23]=g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))));

assign c[24]=g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))));

assign c[25]=g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[26]=g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[27]=g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[28]=g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[29]=g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[30]=g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[31]=g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[32]=g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))); 

assign c[33]=g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[34]=g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[35]=g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[36]=g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[37]=g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[38]=g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[39]=g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[40]=g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[41]=g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[42]=g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[43]=g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[44]=g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[45]=g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[46]=g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[47]=g[47]|(p[47]&(g[46]|(p[46]&(g[45]|(p[45]&(g[44]|(p[44]&(g[43]|(p[43]&(g[42]|(p[42]&(g[41]|(p[41]&(g[40]|(p[40]&(g[39]|(p[39]&(g[38]|(p[38]&(g[37]|(p[37]&(g[36]|(p[36]&(g[35]|(p[35]&(g[34]|(p[34]&(g[33]|(p[33]&(g[32]|(p[32]&(g[31]|(p[31]&(g[30]|(p[30]&(g[29]|(p[29]&(g[28]|(p[28]&(g[27]|(p[27]&(g[26]|(p[26]&(g[25]|(p[25]&(g[24]|(p[24]&(g[23]|(p[23]&(g[22]|(p[22]&(g[21]|(p[21]&(g[20]|(p[20]&(g[19]|(p[19]&(g[18]|(p[18]&(g[17]|(p[17]&(g[16]|(p[16]&(g[15]|(p[15]&(g[14]|(p[14]&(g[13]|(p[13]&(g[12]|(p[12]&(g[11]|(p[11]&(g[10]|(p[10]&(g[9]|(p[9]&(g[8]|(p[8]&(g[7]|(p[7]&(g[6]|(p[6]&(g[5]|(p[5]&(g[4]|(p[4]&(g[3]|(p[3]&(g[2]|(p[2]&(g[1]|(p[1]&(g[0]|(p[0]&cin)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

assign c[48]=cin;

endmodule   

module msum_calculation(p,c,sum);

  output [48:0]sum;

  input [47:0]p;

  input [48:0]c;


  assign sum[0]=p[0]^c[48];

  assign sum[1]=p[1]^c[0];

  assign sum[2]=p[2]^c[1];

  assign sum[3]=p[3]^c[2];

  assign sum[4]=p[4]^c[3];

  assign sum[5]=p[5]^c[4];

  assign sum[6]=p[6]^c[5];

  assign sum[7]=p[7]^c[6];

  assign sum[8]=p[8]^c[7];

  assign sum[9]=p[9]^c[8];

  assign sum[10]=p[10]^c[9];

  assign sum[11]=p[11]^c[10];

  assign sum[12]=p[12]^c[11];

  assign sum[13]=p[13]^c[12];

  assign sum[14]=p[14]^c[13];

  assign sum[15]=p[15]^c[14];

  assign sum[16]=p[16]^c[15];

  assign sum[17]=p[17]^c[16];

  assign sum[18]=p[18]^c[17];

  assign sum[19]=p[19]^c[18];

  assign sum[20]=p[20]^c[19];

  assign sum[21]=p[21]^c[20];

  assign sum[22]=p[22]^c[21];

  assign sum[23]=p[23]^c[22];

  assign sum[24]=p[24]^c[23];

  assign sum[25]=p[25]^c[24];

  assign sum[26]=p[26]^c[25];

  assign sum[27]=p[27]^c[26];

  assign sum[28]=p[28]^c[27];

  assign sum[29]=p[29]^c[28];

  assign sum[30]=p[30]^c[29];

  assign sum[31]=p[31]^c[30];

  assign sum[32]=p[32]^c[31];

  assign sum[33]=p[33]^c[32];

  assign sum[34]=p[34]^c[33];

  assign sum[35]=p[35]^c[34];

  assign sum[36]=p[36]^c[35];

  assign sum[37]=p[37]^c[36];

  assign sum[38]=p[38]^c[37];

  assign sum[39]=p[39]^c[38];

  assign sum[40]=p[40]^c[39];

  assign sum[41]=p[41]^c[40];

  assign sum[42]=p[42]^c[41];

  assign sum[43]=p[43]^c[42];

  assign sum[44]=p[44]^c[43];

  assign sum[45]=p[45]^c[44];

  assign sum[46]=p[46]^c[45];

  assign sum[47]=p[47]^c[46];


  assign sum[48]=c[47];

endmodule

module mcla64(a,b,cin,sum);

  input [47:0]a,b;

  input cin;

  output [48:0]sum;

  wire [47:0]p;

  wire [48:0]c;
   

mcarry_calculation cc(a,b,p,cin,c);  

msum_calculation sc(p,c,sum);  
  
endmodule

module mfulladder(a,b,cin,s,cout);

input a,b,cin;

output s,cout;

assign s=a^b^cin;

assign cout=(a&b)|(b&cin)|(cin&a);

endmodule


module mcsaveadder(X,Y,Z,U,V);

input [47:0]X;

input [47:0]Y;

input [47:0]Z;

output [47:0]U;

output [47:0]V;

wire m;

assign V[0] = 0;

mfulladder fa0(X[0],Y[0],Z[0],U[0],V[1]);

mfulladder fa1(X[1],Y[1],Z[1],U[1],V[2]);

mfulladder fa2(X[2],Y[2],Z[2],U[2],V[3]);

mfulladder fa3(X[3],Y[3],Z[3],U[3],V[4]);

mfulladder fa4(X[4],Y[4],Z[4],U[4],V[5]);

mfulladder fa5(X[5],Y[5],Z[5],U[5],V[6]);

mfulladder fa6(X[6],Y[6],Z[6],U[6],V[7]);

mfulladder fa7(X[7],Y[7],Z[7],U[7],V[8]);

mfulladder fa8(X[8],Y[8],Z[8],U[8],V[9]);

mfulladder fa9(X[9],Y[9],Z[9],U[9],V[10]);

mfulladder fa10(X[10],Y[10],Z[10],U[10],V[11]);

mfulladder fa11(X[11],Y[11],Z[11],U[11],V[12]);

mfulladder fa12(X[12],Y[12],Z[12],U[12],V[13]);

mfulladder fa13(X[13],Y[13],Z[13],U[13],V[14]);

mfulladder fa14(X[14],Y[14],Z[14],U[14],V[15]);

mfulladder fa15(X[15],Y[15],Z[15],U[15],V[16]);

mfulladder fa16(X[16],Y[16],Z[16],U[16],V[17]);

mfulladder fa17(X[17],Y[17],Z[17],U[17],V[18]);

mfulladder fa18(X[18],Y[18],Z[18],U[18],V[19]);

mfulladder fa19(X[19],Y[19],Z[19],U[19],V[20]);

mfulladder fa20(X[20],Y[20],Z[20],U[20],V[21]);

mfulladder fa21(X[21],Y[21],Z[21],U[21],V[22]);

mfulladder fa22(X[22],Y[22],Z[22],U[22],V[23]);

mfulladder fa23(X[23],Y[23],Z[23],U[23],V[24]);

mfulladder fa24(X[24],Y[24],Z[24],U[24],V[25]);

mfulladder fa25(X[25],Y[25],Z[25],U[25],V[26]);

mfulladder fa26(X[26],Y[26],Z[26],U[26],V[27]);

mfulladder fa27(X[27],Y[27],Z[27],U[27],V[28]);

mfulladder fa28(X[28],Y[28],Z[28],U[28],V[29]);

mfulladder fa29(X[29],Y[29],Z[29],U[29],V[30]);

mfulladder fa30(X[30],Y[30],Z[30],U[30],V[31]);

mfulladder fa31(X[31],Y[31],Z[31],U[31],V[32]);

mfulladder fa32(X[32],Y[32],Z[32],U[32],V[33]);

mfulladder fa33(X[33],Y[33],Z[33],U[33],V[34]);

mfulladder fa34(X[34],Y[34],Z[34],U[34],V[35]);

mfulladder fa35(X[35],Y[35],Z[35],U[35],V[36]);

mfulladder fa36(X[36],Y[36],Z[36],U[36],V[37]);

mfulladder fa37(X[37],Y[37],Z[37],U[37],V[38]);

mfulladder fa38(X[38],Y[38],Z[38],U[38],V[39]);

mfulladder fa39(X[39],Y[39],Z[39],U[39],V[40]);

mfulladder fa40(X[40],Y[40],Z[40],U[40],V[41]);

mfulladder fa41(X[41],Y[41],Z[41],U[41],V[42]);

mfulladder fa42(X[42],Y[42],Z[42],U[42],V[43]);

mfulladder fa43(X[43],Y[43],Z[43],U[43],V[44]);

mfulladder fa44(X[44],Y[44],Z[44],U[44],V[45]);

mfulladder fa45(X[45],Y[45],Z[45],U[45],V[46]);

mfulladder fa46(X[46],Y[46],Z[46],U[46],V[47]);

mfulladder fa47(X[47],Y[47],Z[47],U[47],m);

endmodule


module mpartial_product_add(P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23,U0,U1,U2,U3,U4,U5,U6,U7,U8,U9,U10,U11,U12,U13,U14,U15,U16,U17,U18,U19,U20,U29,V0,V1,V2,V3,V4,V5,V6,V7,V8,V9,V10,V11,V12,V13,V14,V15,V16,V17,V18,V19,V20,V29);

input [47:0]P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23;

output [47:0]U0,U1,U2,U3,U4,U5,U6,U7,U8,U9,U10,U11,U12,U13,U14,U15,U16,U17,U18,U19,U20,U29;

output [47:0]V0,V1,V2,V3,V4,V5,V6,V7,V8,V9,V10,V11,V12,V13,V14,V15,V16,V17,V18,V19,V20,V29;

mcsaveadder c1(P0,P1,P2,U0,V0);
mcsaveadder c2(P3,P4,P5,U1,V1);
mcsaveadder c3(P6,P7,P8,U2,V2);
mcsaveadder c4(P9,P10,P11,U3,V3);
mcsaveadder c5(P12,P13,P14,U4,V4);
mcsaveadder c6(P15,P16,P17,U5,V5);
mcsaveadder c7(P18,P19,P20,U6,V6);
mcsaveadder c8(P21,P22,P23,U7,V7);

mcsaveadder c9(U0,V0,U1,U8,V8);
mcsaveadder c10(V1,U2,V2,U9,V9);
mcsaveadder c11(U3,V3,U4,U10,V10);
mcsaveadder c12(V4,U5,V5,U11,V11);
mcsaveadder c13(U6,V6,U7,U12,V12);


mcsaveadder c14(U8,V8,U9,U13,V13);
mcsaveadder c15(V9,U10,V10,U14,V14);
mcsaveadder c16(U11,V11,U12,U15,V15);

mcsaveadder c17(U13,V13,U14,U16,V16);
mcsaveadder c18(V14,U15,V15,U17,V17);


mcsaveadder c19(U16,V16,U17,U18,V18);
mcsaveadder c20(V17,V12,V7,U19,V19);

mcsaveadder c21(U18,V18,U19,U20,V20);

mcsaveadder c22(U20,V20,V19,U29,V29);


endmodule


module mpartial_product_gen(A,B,P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23);

output [47:0]P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23;

input [23:0]A,B;

assign P0=B[0]?A:48'd0;
																																																																																																																																			
assign P1=B[1]?A<<1:48'd0;

assign P2=B[2]?A<<2:48'd0;

assign P3=B[3]?A<<3:48'd0;

assign P4=B[4]?A<<4:48'd0;

assign P5=B[5]?A<<5:48'd0;

assign P6=B[6]?A<<6:48'd0;

assign P7=B[7]?A<<7:48'd0;

assign P8=B[8]?A<<8:48'd0;

assign P9=B[9]?A<<9:48'd0;

assign P10=B[10]?A<<10:48'd0;

assign P11=B[11]?A<<11:48'd0;

assign P12=B[12]?A<<12:48'd0;

assign P13=B[13]?A<<13:48'd0;

assign P14=B[14]?A<<14:48'd0;

assign P15=B[15]?A<<15:48'd0;

assign P16=B[16]?A<<16:48'd0;

assign P17=B[17]?A<<17:48'd0;

assign P18=B[18]?A<<18:48'd0;

assign P19=B[19]?A<<19:48'd0;

assign P20=B[20]?A<<20:48'd0;

assign P21=B[21]?A<<21:48'd0;

assign P22=B[22]?A<<22:48'd0;

assign P23=B[23]?A<<23:48'd0;

endmodule


module mwallace_tree_mult32(A,B,product);

input [23:0]A,B;

wire [47:0]U0,U1,U2,U3,U4,U5,U6,U7,U8,U9,U10,U11,U12,U13,U14,U15,U16,U17,U18,U19,U20,U29;

wire [47:0]V0,V1,V2,V3,V4,V5,V6,V7,V8,V9,V10,V11,V12,V13,V14,V15,V16,V17,V18,V19,V20,V29;

wire carry_wire;

wire [48:0]product_wire;

reg [47:0]product_reg;

reg carry_reg;

output [48:0]product;

wire carry;

wire [47:0]P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23;

reg [47:0]regU29,regV29;


mpartial_product_gen ppgen(A,B,P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23);

mpartial_product_add ppadd(P0,P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16,P17,P18,P19,P20,P21,P22,P23,U0,U1,U2,U3,U4,U5,U6,U7,U8,U9,U10,U11,U12,U13,U14,U15,U16,U17,U18,U19,U20,U29,V0,V1,V2,V3,V4,V5,V6,V7,V8,V9,V10,V11,V12,V13,V14,V15,V16,V17,V18,V19,V20,V29);

mcla64 cla(U29,V29,0,product_wire);

assign product=product_wire;

endmodule


module madd(Sa,Sb,Sc,MaOut,MbOut,Mc);
input Sa,Sb;
output reg Sc;   
input [23:0]MaOut,MbOut;
reg [23:0]M1,M2;
wire [48:0]M;
output reg [48:0]Mc;
wire sin;
assign sin = Sa^Sb;

always@ (*)
begin
	//$display("sin=%b\n",sin);
	if(sin)
	begin
		M1=MaOut;
	   	M2=MbOut;
	    Mc=M;
	    Sc=1'b1;	
		
	end
	
	else
	begin
	   	M1=MaOut;
		M2=MbOut; 
		Mc=M;
		Sc=1'b0;
	end
end

mwallace_tree_mult32 wc(M1,M2,M);	

endmodule

module exponent_add(Sa,Sb,SaOut,SbOut,Ma,Mb,Ea,Eb,Ec,MaOut,MbOut);
input Sa,Sb;
output SaOut,SbOut;
input [23:0]Ma,Mb;
output [23:0]MaOut,MbOut;
input [7:0]Ea,Eb;
wire [7:0]EaOut,EbOut;
output [7:0]Ec;

assign EaOut = Ea-8'b11111111;
assign EbOut = Eb-8'b11111111;
assign Ec = EaOut+EbOut+8'b11111111;
assign MaOut = Ma;
assign MbOut = Mb;
assign SaOut = Sa;
assign SbOut = Sb;

endmodule        

module fpm(a,b,c);
input [31:0]a,b;
input clk;
output [31:0]c;
wire [31:0]cwire;
reg [31:0]cReg;
wire Sa,Sb,Sc;
wire [7:0]Ea,Eb,Ec;
wire [23:0]Ma,Mb,MaOut,MbOut;
wire [48:0]Mc;
wire [24:0]Mc1;
reg [24:0]Mc1Reg;
reg [48:0]McReg;
reg ScReg;
//wire s;
wire [48:0]McOut;
wire [7:0]EcOut;
wire ScOut,SaOut,SbOut;
reg SaOutReg,SbOutReg,ScOutReg;
reg [7:0]EcReg,EcReg1,EcOutReg;
reg [23:0]MaOutReg,MbOutReg;
assign Ma[23]=1'b1;
assign Mb[23]=1'b1;
assign Sa=a[31];
assign Sb=b[31];
assign Ma[22:0]=a[22:0];
assign Mb[22:0]=b[22:0];
assign Ea=a[30:23];
assign Eb=b[30:23];

exponent_add cs(Sa,Sb,SaOut,SbOut,Ma,Mb,Ea,Eb,Ec,MaOut,MbOut);

madd ad(SaOutReg,SbOutReg,Sc,MaOutReg,MbOutReg,Mc);

mresult_normalize rn(McReg,ScReg,EcReg1,ScOut,EcOut,Mc1);

//combine cp(ScOutReg,EcOutReg,Mc1Reg,cwire);
assign c={ScOutReg,EcOutReg,Mc1Reg[22:0]};

always @(*)
begin
	//stage 1
	 SaOutReg<=SaOut;
	 SbOutReg<=SbOut;
	 MaOutReg<=MaOut;
	 MbOutReg<=MbOut;
	 EcReg<=Ec;

	 //stage 2
	 ScReg<=Sc;
	 McReg<=Mc;
	 EcReg1<=EcReg;

	 //stage3
	 ScOutReg<=ScOut;
	 EcOutReg<=EcOut;
	 Mc1Reg<=Mc1;

	 //stage4
	

end

endmodule       






































